
module output_lut(din, clk, rst, ena, dout);
    parameter NDATA = 128;
    parameter NDATA_LOG = $clog2(NDATA);

    input [NDATA_LOG-1:0] din;
    input clk;
    input rst;
    input ena;

    output reg [8:0] dout = 9'd0;

    always @ (posedge clk or negedge rst) begin
        if (!rst)
            dout <= 9'd0;
        else
            if (!ena)
                case (din)
                    0: dout <= 9'd90;
                    1: dout <= 9'd89;
                    2: dout <= 9'd88;
                    3: dout <= 9'd87;
                    4: dout <= 9'd86;
                    5: dout <= 9'd85;
                    6: dout <= 9'd85;
                    7: dout <= 9'd84;
                    8: dout <= 9'd83;
                    9: dout <= 9'd82;
                    10: dout <= 9'd81;
                    11: dout <= 9'd80;
                    12: dout <= 9'd79;
                    13: dout <= 9'd78;
                    14: dout <= 9'd77;
                    15: dout <= 9'd76;
                    16: dout <= 9'd75;
                    17: dout <= 9'd74;
                    18: dout <= 9'd73;
                    19: dout <= 9'd72;
                    20: dout <= 9'd71;
                    21: dout <= 9'd71;
                    22: dout <= 9'd70;
                    23: dout <= 9'd69;
                    24: dout <= 9'd68;
                    25: dout <= 9'd67;
                    26: dout <= 9'd66;
                    27: dout <= 9'd65;
                    28: dout <= 9'd64;
                    29: dout <= 9'd63;
                    30: dout <= 9'd62;
                    31: dout <= 9'd61;
                    32: dout <= 9'd59;
                    33: dout <= 9'd58;
                    34: dout <= 9'd57;
                    35: dout <= 9'd56;
                    36: dout <= 9'd55;
                    37: dout <= 9'd54;
                    38: dout <= 9'd53;
                    39: dout <= 9'd52;
                    40: dout <= 9'd51;
                    41: dout <= 9'd49;
                    42: dout <= 9'd48;
                    43: dout <= 9'd47;
                    44: dout <= 9'd46;
                    45: dout <= 9'd44;
                    46: dout <= 9'd43;
                    47: dout <= 9'd42;
                    48: dout <= 9'd40;
                    49: dout <= 9'd39;
                    50: dout <= 9'd37;
                    51: dout <= 9'd36;
                    52: dout <= 9'd34;
                    53: dout <= 9'd33;
                    54: dout <= 9'd31;
                    55: dout <= 9'd29;
                    56: dout <= 9'd27;
                    57: dout <= 9'd25;
                    58: dout <= 9'd23;
                    59: dout <= 9'd21;
                    60: dout <= 9'd18;
                    61: dout <= 9'd14;
                    62: dout <= 9'd10;
                    63: dout <= 9'd0;
                    64: dout <= 9'd0;
                    65: dout <= 9'd180;
                    66: dout <= 9'd170;
                    67: dout <= 9'd166;
                    68: dout <= 9'd162;
                    69: dout <= 9'd159;
                    70: dout <= 9'd157;
                    71: dout <= 9'd155;
                    72: dout <= 9'd153;
                    73: dout <= 9'd151;
                    74: dout <= 9'd149;
                    75: dout <= 9'd147;
                    76: dout <= 9'd146;
                    77: dout <= 9'd144;
                    78: dout <= 9'd143;
                    79: dout <= 9'd141;
                    80: dout <= 9'd140;
                    81: dout <= 9'd138;
                    82: dout <= 9'd137;
                    83: dout <= 9'd136;
                    84: dout <= 9'd134;
                    85: dout <= 9'd133;
                    86: dout <= 9'd132;
                    87: dout <= 9'd131;
                    88: dout <= 9'd129;
                    89: dout <= 9'd128;
                    90: dout <= 9'd127;
                    91: dout <= 9'd126;
                    92: dout <= 9'd125;
                    93: dout <= 9'd124;
                    94: dout <= 9'd123;
                    95: dout <= 9'd122;
                    96: dout <= 9'd121;
                    97: dout <= 9'd119;
                    98: dout <= 9'd118;
                    99: dout <= 9'd117;
                    100: dout <= 9'd116;
                    101: dout <= 9'd115;
                    102: dout <= 9'd114;
                    103: dout <= 9'd113;
                    104: dout <= 9'd112;
                    105: dout <= 9'd111;
                    106: dout <= 9'd110;
                    107: dout <= 9'd109;
                    108: dout <= 9'd109;
                    109: dout <= 9'd108;
                    110: dout <= 9'd107;
                    111: dout <= 9'd106;
                    112: dout <= 9'd105;
                    113: dout <= 9'd104;
                    114: dout <= 9'd103;
                    115: dout <= 9'd102;
                    116: dout <= 9'd101;
                    117: dout <= 9'd100;
                    118: dout <= 9'd99;
                    119: dout <= 9'd98;
                    120: dout <= 9'd97;
                    121: dout <= 9'd96;
                    122: dout <= 9'd95;
                    123: dout <= 9'd95;
                    124: dout <= 9'd94;
                    125: dout <= 9'd93;
                    126: dout <= 9'd92;
                    127: dout <= 9'd91;
                endcase
    end

endmodule
