/**
 *  Electronics Design Competition 2015
 *  Sound Source Localization
 *
 *  Top Level Design: ssl.v
 *  @brief  This module contains the top level design that will be implemented
 *          the FPGA board.
 */

`timescale 1ns/100ps

module ssl(clk, rst, ena);
    input clk;
    input rst;
    input ena;
    

endmodule
